`include "sprot_rand_seq.sv"
