/* 
* Copyright (c) 2004-2023 CVC, VerifWorks, London-UK & Bangalore, India
* http://www.verifworks.com 
* Contact: support@verifworks.com 
* 
* This program is part of Go2UVM at https://github.com/go2uvm/go2uvm
* Some portions of Go2UVM are free software.
* You can redistribute it and/or modify  
* it under the terms of the GNU Lesser General Public License as   
* published by the Free Software Foundation, version 3.
*
* VerifWorks reserves the right to obfuscate part or full of the code
* at any point in time. 
* We also support a comemrical licensing option for an enhanced version
* of Go2UVM, please contact us via support@verifworks.com

* This program is distributed in the hope that it will be useful, but 
* WITHOUT ANY WARRANTY; without even the implied warranty of 
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU 
* Lesser General Lesser Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program. If not, see <http://www.gnu.org/licenses/>.
*/


import apb2_master_pkg::*;
interface apb2_master_if (input logic pclk);
 
  logic pselx;
  logic presetn;
  logic pwrite;
  logic penable;
  logic [DATA_WIDTH-1:0] pwdata;
  logic [ADDR_WIDTH-1:0] paddr;
  logic [DATA_WIDTH-1:0] prdata;

//Clocking block declaration
  clocking apb_driver_cb @(posedge pclk);
    output presetn;
    output pwrite;
    output penable;
    output pwdata;
    output paddr;
    output pselx;
    input prdata;
  endclocking:apb_driver_cb

  clocking apb_monitor_cb @(posedge pclk);
    input presetn;
    input pwrite;
    input penable;
    input pwdata;
    input paddr;
    input pselx;
    input prdata;
  endclocking:apb_monitor_cb 

endinterface : apb2_master_if
