// Copyright (c) 2004-2017 VerifWorks, Bangalore, India
// http://www.verifworks.com 
// Contact: support@verifworks.com 
// 
// This program is part of Go2UVM at www.go2uvm.org
// Some portions of Go2UVM are free software.
// You can redistribute it and/or modify  
// it under the terms of the GNU Lesser General Public License as   
// published by the Free Software Foundation, version 3.
//
// VerifWorks reserves the right to obfuscate part or full of the code
// at any point in time. 
// We also support a comemrical licensing option for an enhanced version
// of Go2UVM, please contact us via support@verifworks.com
//
// This program is distributed in the hope that it will be useful, but 
// WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU 
// Lesser General Lesser Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public License
// along with this program. If not, see <http://www.gnu.org/licenses/>.

/********************************************
* VerifWorks Go2UVM App: VW_DVC_Go2UVM
* Automatically generated by VerifWorks's DVC_Go2UVM Riviera Apps 
* Thanks for using VerifWorks products
* Visit http://www.verifworks.com for more 
* Generated on   : 2016-06-21 21:50:32
********************************************/ 


// Generating Go2UVM Test for module: sprot
// ---------------------------------------------------------

// Automatically generated from VerifWorks's DVCreate-Go2UVM product
// Thanks for using VerifWorks products, see http://www.verifworks.com for more

import uvm_pkg::*;
`include "vw_go2uvm_macros.svh"
// Import Go2UVM Package
import vw_go2uvm_pkg::*;

// Use the base class provided by the vw_go2uvm_pkg
`G2U_TEST_BEGIN(sprot_test)
  // Create a handle to the actual interface
   `G2U_GET_VIF(sprot_if)
   
  logic [7:0] local_byte_val;

  task reset;
    `g2u_display ("Start of reset")
     this.vif.cb.rst_n <= 1'b0;
     repeat (5) @ (this.vif.cb);
     this.vif.cb.rst_n <= 1'b1;
     repeat (1) @ (this.vif.cb);
    `g2u_display ("End of reset")
  endtask : reset

  task main ();
    `g2u_display("Starting force test");
    g2u_force("sprot_go2uvm.aldec_src_ex", 22);
    g2u_force("sprot_go2uvm.sprot_0.byte_val", 22);
    #100;
    g2u_force("sprot_go2uvm.sprot_0.byte_val", 'haa);
    #100;
    `g2u_display ("End of main")
  endtask : main
   
`G2U_TEST_END

