/*
This file is not part of current release of Go2UVM. We do have a limited customer availability of this feature, please contact support@verifworks.com for more details


*/
