//#----------------------------------------------------------------------
//#   Copyright 2004-2014 CVC Pvt. Ltd. Bangalore, India
//#    http://www.cvcblr.com 
//#   All Rights Reserved Worldwide
//#
//#   Licensed under the Apache License, Version 2.0 (the
//#   "License"); you may not use this file except in
//#   compliance with the License.  You may obtain a copy of
//#   the License at
//#
//#       http://www.apache.org/licenses/LICENSE-2.0
//#
//#   Unless required by applicable law or agreed to in
//#   writing, software distributed under the License is
//#   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//#   CONDITIONS OF ANY KIND, either express or implied.  See
//#   the License for the specific language governing
//#   permissions and limitations under the License.
//#----------------------------------------------------------------------

`include "sprot_xactn.sv"
`include "sprot_sequencer.sv"
`include "sprot_input_monitor.sv"
`include "sprot_output_monitor.sv"
`include "sprot_fcov.sv"
`include "sprot_scoreboard.sv"
`include "sprot_driver.sv"
`include "sprot_agent.sv"
`include "sprot_env.sv"
`include "sprot_seq_lib.sv"
`include "sprot_base_test.sv"
