/* 
* Copyright (c) 2004-2017 VerifWorks, Bangalore, India
* http://www.verifworks.com 
* Contact: support@verifworks.com 
* 
* This program is part of Go2UVM at www.go2uvm.org
* Some portions of Go2UVM are free software.
* You can redistribute it and/or modify  
* it under the terms of the GNU Lesser General Public License as   
* published by the Free Software Foundation, version 3.
*
* VerifWorks reserves the right to obfuscate part or full of the code
* at any point in time. 
* We also support a comemrical licensing option for an enhanced version
* of Go2UVM, please contact us via support@verifworks.com

* This program is distributed in the hope that it will be useful, but 
* WITHOUT ANY WARRANTY; without even the implied warranty of 
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU 
* Lesser General Lesser Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program. If not, see <http://www.gnu.org/licenses/>.
*/


//---------------------------------------------------------------------------
//   THIS IS AN AUTOMATICALLY GENERATED CODE
//   Generated by GenReg, a product from VerifWorks http://www.verifworks.com
//   A venture of CVC Pvt. Ltd. http://www.cvcblr.com
//   UVM Register Kit Version 1.1
//---------------------------------------------------------------------------
// Project           : i2c_spec_reg_model
// Unit              : i2c_spec_pkg_uvm
// File              : i2c_spec_reg_model
// Created by        : student
// Date of creation  : 7/19/2105 4:12 PM
//--------------------------------------------------------------------------- 
// Title             : cvc_reg_model
//
// Description       : 
//
//---------------------------------------------------------------------------

//---------------------------------------------------------------------------
//i2c_spec_pkg_uvm
//---------------------------------------------------------------------------

   import uvm_pkg::*;

   `include "uvm_macros.svh"

   /* DEFINE REGISTER CLASSES */
   //---------------------------------------------------------------------------
   // Class: i2c_spec_PRERlo_reg
   //---------------------------------------------------------------------------

   class i2c_spec_PRERlo_reg extends uvm_reg;
      `uvm_object_utils (i2c_spec_PRERlo_reg)

      rand uvm_reg_field Prescale_register;


      // Function: new
      //
      function new(string name = "i2c_spec_PRERlo_reg");
         super.new(name,8,UVM_NO_COVERAGE);
      endfunction : new


      // Function: build
      //
      virtual function void build();

         this.Prescale_register = uvm_reg_field::type_id::create("Prescale_register");

         Prescale_register.configure(.parent(this),.size(8),.lsb_pos(0),.access("RW"),.volatile(0),.reset(8'hff),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
      endfunction : build
   endclass



   //---------------------------------------------------------------------------
   // Class: i2c_spec_PRERhi_reg
   //---------------------------------------------------------------------------

   class i2c_spec_PRERhi_reg extends uvm_reg;
      `uvm_object_utils (i2c_spec_PRERhi_reg)

      rand uvm_reg_field Prescale_register;


      // Function: new
      //
      function new(string name = "i2c_spec_PRERhi_reg");
         super.new(name,8,UVM_NO_COVERAGE);
      endfunction : new


      // Function: build
      //
      virtual function void build();

         this.Prescale_register = uvm_reg_field::type_id::create("Prescale_register");

         Prescale_register.configure(.parent(this),.size(8),.lsb_pos(0),.access("RW"),.volatile(0),.reset(8'hff),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
      endfunction : build
   endclass



   //---------------------------------------------------------------------------
   // Class: i2c_spec_CTR_reg
   //---------------------------------------------------------------------------

   class i2c_spec_CTR_reg extends uvm_reg;
      `uvm_object_utils (i2c_spec_CTR_reg)

      rand uvm_reg_field EN;
      rand uvm_reg_field IEN;
      rand uvm_reg_field Reserved;


      // Function: new
      //
      function new(string name = "i2c_spec_CTR_reg");
         super.new(name,8,UVM_NO_COVERAGE);
      endfunction : new


      // Function: build
      //
      virtual function void build();

         this.EN = uvm_reg_field::type_id::create("EN");
         this.IEN = uvm_reg_field::type_id::create("IEN");
         this.Reserved = uvm_reg_field::type_id::create("Reserved");

         EN.configure(.parent(this),.size(1),.lsb_pos(7),.access("RW"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
         IEN.configure(.parent(this),.size(1),.lsb_pos(6),.access("RW"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
         Reserved.configure(.parent(this),.size(6),.lsb_pos(0),.access("RW"),.volatile(0),.reset(6'b000000),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
      endfunction : build
   endclass



   //---------------------------------------------------------------------------
   // Class: i2c_spec_TXR_reg
   //---------------------------------------------------------------------------

   class i2c_spec_TXR_reg extends uvm_reg;
      `uvm_object_utils (i2c_spec_TXR_reg)

      rand uvm_reg_field Transmit_register_0;
      rand uvm_reg_field Transmit_register_1;


      // Function: new
      //
      function new(string name = "i2c_spec_TXR_reg");
         super.new(name,8,UVM_NO_COVERAGE);
      endfunction : new


      // Function: build
      //
      virtual function void build();

         this.Transmit_register_0 = uvm_reg_field::type_id::create("Transmit_register_0");
         this.Transmit_register_1 = uvm_reg_field::type_id::create("Transmit_register_1");

         Transmit_register_0.configure(.parent(this),.size(7),.lsb_pos(1),.access("WO"),.volatile(0),.reset(7'b0000000),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
         Transmit_register_1.configure(.parent(this),.size(1),.lsb_pos(0),.access("WO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
      endfunction : build
   endclass



   //---------------------------------------------------------------------------
   // Class: i2c_spec_RXR_reg
   //---------------------------------------------------------------------------

   class i2c_spec_RXR_reg extends uvm_reg;
      `uvm_object_utils (i2c_spec_RXR_reg)

           uvm_reg_field Receive_register;


      // Function: new
      //
      function new(string name = "i2c_spec_RXR_reg");
         super.new(name,8,UVM_NO_COVERAGE);
      endfunction : new


      // Function: build
      //
      virtual function void build();

         this.Receive_register = uvm_reg_field::type_id::create("Receive_register");

         Receive_register.configure(.parent(this),.size(8),.lsb_pos(0),.access("RO"),.volatile(0),.reset(8'h00),.has_reset(0),.is_rand(0),
                      .individually_accessible(0)); 
      endfunction : build
   endclass



   //---------------------------------------------------------------------------
   // Class: i2c_spec_CR_reg
   //---------------------------------------------------------------------------

   class i2c_spec_CR_reg extends uvm_reg;
      `uvm_object_utils (i2c_spec_CR_reg)

      rand uvm_reg_field STA;
      rand uvm_reg_field STO;
      rand uvm_reg_field RD;
      rand uvm_reg_field WR;
      rand uvm_reg_field ACK;
      rand uvm_reg_field Reserved;
      rand uvm_reg_field IACK;


      // Function: new
      //
      function new(string name = "i2c_spec_CR_reg");
         super.new(name,8,UVM_NO_COVERAGE);
      endfunction : new


      // Function: build
      //
      virtual function void build();

         this.STA = uvm_reg_field::type_id::create("STA");
         this.STO = uvm_reg_field::type_id::create("STO");
         this.RD = uvm_reg_field::type_id::create("RD");
         this.WR = uvm_reg_field::type_id::create("WR");
         this.ACK = uvm_reg_field::type_id::create("ACK");
         this.Reserved = uvm_reg_field::type_id::create("Reserved");
         this.IACK = uvm_reg_field::type_id::create("IACK");

         STA.configure(.parent(this),.size(1),.lsb_pos(7),.access("WO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
         STO.configure(.parent(this),.size(1),.lsb_pos(6),.access("WO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
         RD.configure(.parent(this),.size(1),.lsb_pos(5),.access("WO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
         WR.configure(.parent(this),.size(1),.lsb_pos(4),.access("WO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
         ACK.configure(.parent(this),.size(1),.lsb_pos(3),.access("WO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
         Reserved.configure(.parent(this),.size(2),.lsb_pos(1),.access("WO"),.volatile(0),.reset(2'b00),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
         IACK.configure(.parent(this),.size(1),.lsb_pos(0),.access("WO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(1),
                      .individually_accessible(0)); 
      endfunction : build
   endclass



   //---------------------------------------------------------------------------
   // Class: i2c_spec_SR_reg
   //---------------------------------------------------------------------------

   class i2c_spec_SR_reg extends uvm_reg;
      `uvm_object_utils (i2c_spec_SR_reg)

           uvm_reg_field RxACK;
           uvm_reg_field Busy;
           uvm_reg_field AL;
           uvm_reg_field Reserved;
           uvm_reg_field TIP;
           uvm_reg_field I_F;


      // Function: new
      //
      function new(string name = "i2c_spec_SR_reg");
         super.new(name,8,UVM_NO_COVERAGE);
      endfunction : new


      // Function: build
      //
      virtual function void build();

         this.RxACK = uvm_reg_field::type_id::create("RxACK");
         this.Busy = uvm_reg_field::type_id::create("Busy");
         this.AL = uvm_reg_field::type_id::create("AL");
         this.Reserved = uvm_reg_field::type_id::create("Reserved");
         this.TIP = uvm_reg_field::type_id::create("TIP");
         this.I_F = uvm_reg_field::type_id::create("I_F");

         RxACK.configure(.parent(this),.size(1),.lsb_pos(7),.access("RO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(0),
                      .individually_accessible(0)); 
         Busy.configure(.parent(this),.size(1),.lsb_pos(6),.access("RO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(0),
                      .individually_accessible(0)); 
         AL.configure(.parent(this),.size(1),.lsb_pos(5),.access("RO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(0),
                      .individually_accessible(0)); 
         Reserved.configure(.parent(this),.size(3),.lsb_pos(2),.access("RO"),.volatile(0),.reset(3'b000),.has_reset(0),.is_rand(0),
                      .individually_accessible(0)); 
         TIP.configure(.parent(this),.size(1),.lsb_pos(1),.access("RO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(0),
                      .individually_accessible(0)); 
         I_F.configure(.parent(this),.size(1),.lsb_pos(0),.access("RO"),.volatile(0),.reset(1'b0),.has_reset(0),.is_rand(0),
                      .individually_accessible(0)); 
      endfunction : build
   endclass



    /* BLOCKS */

    //----------------------------------------------------------------------
    // Class :i2c_reg_block

    //----------------------------------------------------------------------

   class i2c_reg_block extends uvm_reg_block;
      `uvm_object_utils(i2c_reg_block)

      rand i2c_spec_PRERlo_reg i2c_spec_PRERlo;
      rand i2c_spec_PRERhi_reg i2c_spec_PRERhi;
      rand i2c_spec_CTR_reg i2c_spec_CTR;
      rand i2c_spec_TXR_reg i2c_spec_TXR;
      rand i2c_spec_RXR_reg i2c_spec_RXR;
      rand i2c_spec_CR_reg i2c_spec_CR;
      rand i2c_spec_SR_reg i2c_spec_SR;


      uvm_reg_map i2c_reg_block_map;


      // Function: new
      //
      function new(string name = "i2c_reg_block");
         super.new(name, UVM_NO_COVERAGE);
      endfunction



      // Function: build
      //
      virtual function void build();
         i2c_spec_PRERlo = i2c_spec_PRERlo_reg::type_id::create("i2c_spec_PRERlo");
         i2c_spec_PRERlo.configure(this);
         i2c_spec_PRERlo.build();


         i2c_spec_PRERhi = i2c_spec_PRERhi_reg::type_id::create("i2c_spec_PRERhi");
         i2c_spec_PRERhi.configure(this);
         i2c_spec_PRERhi.build();


         i2c_spec_CTR = i2c_spec_CTR_reg::type_id::create("i2c_spec_CTR");
         i2c_spec_CTR.configure(this);
         i2c_spec_CTR.build();


         i2c_spec_TXR = i2c_spec_TXR_reg::type_id::create("i2c_spec_TXR");
         i2c_spec_TXR.configure(this);
         i2c_spec_TXR.build();


         i2c_spec_RXR = i2c_spec_RXR_reg::type_id::create("i2c_spec_RXR");
         i2c_spec_RXR.configure(this);
         i2c_spec_RXR.build();


         i2c_spec_CR = i2c_spec_CR_reg::type_id::create("i2c_spec_CR");
         i2c_spec_CR.configure(this);
         i2c_spec_CR.build();


         i2c_spec_SR = i2c_spec_SR_reg::type_id::create("i2c_spec_SR");
         i2c_spec_SR.configure(this);
         i2c_spec_SR.build();


         i2c_reg_block_map = create_map("i2c_reg_block_map",'h0,4,UVM_LITTLE_ENDIAN);
         default_map =i2c_reg_block_map;
         i2c_reg_block_map.add_reg(i2c_spec_PRERlo,'h0,"RW");
         i2c_reg_block_map.add_reg(i2c_spec_PRERhi,'h1,"RW");
         i2c_reg_block_map.add_reg(i2c_spec_CTR,'h2,"RW");
         i2c_reg_block_map.add_reg(i2c_spec_TXR,'h3,"WO");
         i2c_reg_block_map.add_reg(i2c_spec_RXR,'h3,"RO");
         i2c_reg_block_map.add_reg(i2c_spec_CR,'h4,"WO");
         i2c_reg_block_map.add_reg(i2c_spec_SR,'h4,"RO");

         lock_model();
      endfunction
   endclass

